
// 0x400000 - 0x400013 -> the memory map for Pattern matching peripheral

module PMP (
    

)



endmodule